magic
tech sky130A
magscale 1 2
timestamp 1712671220
<< metal1 >>
rect 25390 4656 25690 4662
rect 25690 4356 26882 4656
rect 25390 4350 25690 4356
rect 26896 3406 27016 3548
rect 31042 3446 31312 3566
rect 31432 3446 31438 3566
rect 26890 3286 26896 3406
rect 27016 3286 27022 3406
rect 26164 2712 26464 2718
rect 26464 2412 26992 2712
rect 26164 2406 26464 2412
<< via1 >>
rect 25390 4356 25690 4656
rect 31312 3446 31432 3566
rect 26896 3286 27016 3406
rect 26164 2412 26464 2712
<< metal2 >>
rect 24353 4656 24643 4660
rect 24348 4651 25390 4656
rect 24348 4361 24353 4651
rect 24643 4361 25390 4651
rect 24348 4356 25390 4361
rect 25690 4356 25696 4656
rect 24353 4352 24643 4356
rect 31312 3566 31432 3572
rect 26896 3406 27016 3412
rect 31312 3317 31432 3446
rect 26896 3243 27016 3286
rect 26892 3133 26901 3243
rect 27011 3133 27020 3243
rect 31308 3207 31317 3317
rect 31427 3207 31436 3317
rect 31312 3202 31432 3207
rect 26896 3128 27016 3133
rect 25951 2712 26241 2716
rect 25946 2707 26164 2712
rect 25946 2417 25951 2707
rect 25946 2412 26164 2417
rect 26464 2412 26470 2712
rect 25951 2408 26241 2412
<< via2 >>
rect 24353 4361 24643 4651
rect 26901 3133 27011 3243
rect 31317 3207 31427 3317
rect 25951 2417 26164 2707
rect 26164 2417 26241 2707
<< metal3 >>
rect 6811 4656 7109 4661
rect 6810 4655 24648 4656
rect 6810 4357 6811 4655
rect 7109 4651 24648 4655
rect 7109 4361 24353 4651
rect 24643 4361 24648 4651
rect 7109 4357 24648 4361
rect 6810 4356 24648 4357
rect 6811 4351 7109 4356
rect 31312 3317 31432 3322
rect 26896 3243 27016 3248
rect 26896 3133 26901 3243
rect 27011 3133 27016 3243
rect 26896 3021 27016 3133
rect 31312 3207 31317 3317
rect 31427 3207 31432 3317
rect 31312 3097 31432 3207
rect 26891 2903 26897 3021
rect 27015 2903 27021 3021
rect 31312 2979 31313 3097
rect 31431 2979 31432 3097
rect 31312 2978 31432 2979
rect 31313 2973 31431 2978
rect 26896 2902 27016 2903
rect 25719 2712 26017 2717
rect 25718 2711 26246 2712
rect 25718 2413 25719 2711
rect 26017 2707 26246 2711
rect 26241 2417 26246 2707
rect 26017 2413 26246 2417
rect 25718 2412 26246 2413
rect 25719 2407 26017 2412
<< via3 >>
rect 6811 4357 7109 4655
rect 26897 2903 27015 3021
rect 31313 2979 31431 3097
rect 25719 2707 26017 2711
rect 25719 2417 25951 2707
rect 25951 2417 26017 2707
rect 25719 2413 26017 2417
<< metal4 >>
rect 798 44676 858 45152
rect 1534 44676 1594 45152
rect 2270 44676 2330 45152
rect 3006 44676 3066 45152
rect 3742 44676 3802 45152
rect 4478 44676 4538 45152
rect 5214 44676 5274 45152
rect 5950 44676 6010 45152
rect 6686 44676 6746 45152
rect 7422 44676 7482 45152
rect 8158 44676 8218 45152
rect 8894 44676 8954 45152
rect 9630 44676 9690 45152
rect 10366 44676 10426 45152
rect 11102 44676 11162 45152
rect 11838 44676 11898 45152
rect 12574 44676 12634 45152
rect 13310 44676 13370 45152
rect 14046 44676 14106 45152
rect 14782 44676 14842 45152
rect 15518 44676 15578 45152
rect 16254 44676 16314 45152
rect 16990 44676 17050 45152
rect 17726 44676 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 680 44414 17928 44676
rect 200 4656 500 44152
rect 200 4655 7110 4656
rect 200 4357 6811 4655
rect 7109 4357 7110 4655
rect 200 4356 7110 4357
rect 200 1000 500 4356
rect 9800 2712 10100 44414
rect 31312 3097 31432 3098
rect 26896 3021 27016 3022
rect 26896 2903 26897 3021
rect 27015 2903 27016 3021
rect 9800 2711 26018 2712
rect 9800 2413 25719 2711
rect 26017 2413 26018 2711
rect 9800 2412 26018 2413
rect 9800 1000 10100 2412
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 2903
rect 31312 2979 31313 3097
rect 31431 2979 31432 3097
rect 31312 0 31432 2979
use inverter  inverter_0
timestamp 1712074259
transform 1 0 26874 0 1 3208
box -236 -828 4448 1468
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
