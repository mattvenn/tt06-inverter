magic
tech sky130A
magscale 1 2
timestamp 1712320071
<< viali >>
rect 924 964 1044 1008
rect 2108 950 3262 998
rect 930 -370 1040 -328
rect 2134 -386 3270 -334
<< metal1 >>
rect -236 1168 4378 1468
rect 634 798 732 1168
rect 900 1008 1066 1168
rect 1500 1116 1572 1168
rect 1494 1044 1500 1116
rect 1572 1044 1578 1116
rect 2092 1054 3292 1168
rect 900 964 924 1008
rect 1044 964 1066 1008
rect 900 946 1066 964
rect 2090 998 3292 1054
rect 2090 950 2108 998
rect 3262 950 3292 998
rect 2090 944 3292 950
rect 1211 910 1460 911
rect 948 861 1460 910
rect 948 860 1262 861
rect 634 656 962 798
rect 1014 690 1266 770
rect 1346 690 1352 770
rect 720 644 962 656
rect 1411 581 1460 861
rect 951 531 1460 581
rect 1554 855 3749 905
rect 1554 569 1604 855
rect 1762 742 1772 800
rect 1828 742 1838 800
rect 1954 746 1964 804
rect 2020 746 2030 804
rect 2140 744 2150 806
rect 2204 744 2214 806
rect 2342 740 2352 802
rect 2406 740 2416 802
rect 2530 740 2540 802
rect 2594 740 2604 802
rect 2726 744 2736 806
rect 2790 744 2800 806
rect 2910 746 2920 808
rect 2974 746 2984 808
rect 3106 736 3116 798
rect 3170 736 3180 798
rect 3298 740 3308 802
rect 3362 740 3372 802
rect 3490 746 3500 808
rect 3554 746 3564 808
rect 3682 746 3692 808
rect 3746 746 3756 808
rect 1858 620 1868 674
rect 1920 620 1930 674
rect 2050 624 2060 678
rect 2112 624 2122 678
rect 2240 620 2250 674
rect 2302 620 2312 674
rect 2428 616 2438 670
rect 2490 616 2500 670
rect 2624 622 2634 676
rect 2686 622 2696 676
rect 2818 618 2828 672
rect 2880 618 2890 672
rect 3010 614 3020 668
rect 3072 614 3082 668
rect 3206 618 3216 672
rect 3268 618 3278 672
rect 3398 618 3408 672
rect 3460 618 3470 672
rect 3582 618 3592 672
rect 3644 618 3654 672
rect 1543 553 1604 569
rect 76 341 276 392
rect 1347 341 1397 531
rect 1543 503 3663 553
rect 1543 356 1593 503
rect 4142 382 4342 440
rect 76 291 1397 341
rect 76 192 276 291
rect 952 84 1086 90
rect 1347 84 1397 291
rect 1542 350 1622 356
rect 3974 276 4342 382
rect 1542 264 1622 270
rect 1543 84 1593 264
rect 4142 240 4342 276
rect 952 46 1472 84
rect 1042 38 1472 46
rect 1246 34 1472 38
rect 1543 36 3757 84
rect 1543 34 3292 36
rect 3366 34 3757 36
rect 702 -22 954 -2
rect 634 -156 954 -22
rect 1014 -132 1266 -52
rect 1346 -132 1352 -52
rect 634 -528 726 -156
rect 1421 -229 1471 34
rect 1543 -229 1593 34
rect 1756 -64 1766 -6
rect 1822 -64 1832 -6
rect 1948 -60 1958 -2
rect 2014 -60 2024 -2
rect 2134 -62 2144 0
rect 2198 -62 2208 0
rect 2336 -66 2346 -4
rect 2400 -66 2410 -4
rect 2524 -66 2534 -4
rect 2588 -66 2598 -4
rect 2720 -62 2730 0
rect 2784 -62 2794 0
rect 2904 -60 2914 2
rect 2968 -60 2978 2
rect 3100 -70 3110 -8
rect 3164 -70 3174 -8
rect 3292 -66 3302 -4
rect 3356 -66 3366 -4
rect 3484 -60 3494 2
rect 3548 -60 3558 2
rect 3676 -60 3686 2
rect 3740 -60 3750 2
rect 1852 -186 1862 -132
rect 1914 -186 1924 -132
rect 2044 -182 2054 -128
rect 2106 -182 2116 -128
rect 2234 -186 2244 -132
rect 2296 -186 2306 -132
rect 2422 -190 2432 -136
rect 2484 -190 2494 -136
rect 2618 -184 2628 -130
rect 2680 -184 2690 -130
rect 2812 -188 2822 -134
rect 2874 -188 2884 -134
rect 3004 -192 3014 -138
rect 3066 -192 3076 -138
rect 3200 -188 3210 -134
rect 3262 -188 3272 -134
rect 3392 -188 3402 -134
rect 3454 -188 3464 -134
rect 3576 -188 3586 -134
rect 3638 -188 3648 -134
rect 947 -279 1472 -229
rect 1543 -277 3677 -229
rect 1574 -279 3677 -277
rect 908 -328 1060 -320
rect 908 -334 930 -328
rect 906 -370 930 -334
rect 1040 -370 1060 -328
rect 2092 -334 3292 -328
rect 906 -528 1060 -370
rect 1490 -440 1496 -368
rect 1568 -440 1574 -368
rect 2092 -386 2134 -334
rect 3270 -386 3292 -334
rect 1496 -528 1568 -440
rect 2092 -528 3292 -386
rect -166 -828 4448 -528
<< via1 >>
rect 1500 1044 1572 1116
rect 1266 690 1346 770
rect 1772 742 1828 800
rect 1964 746 2020 804
rect 2150 744 2204 806
rect 2352 740 2406 802
rect 2540 740 2594 802
rect 2736 744 2790 806
rect 2920 746 2974 808
rect 3116 736 3170 798
rect 3308 740 3362 802
rect 3500 746 3554 808
rect 3692 746 3746 808
rect 1868 620 1920 674
rect 2060 624 2112 678
rect 2250 620 2302 674
rect 2438 616 2490 670
rect 2634 622 2686 676
rect 2828 618 2880 672
rect 3020 614 3072 668
rect 3216 618 3268 672
rect 3408 618 3460 672
rect 3592 618 3644 672
rect 1542 270 1622 350
rect 1266 -132 1346 -52
rect 1766 -64 1822 -6
rect 1958 -60 2014 -2
rect 2144 -62 2198 0
rect 2346 -66 2400 -4
rect 2534 -66 2588 -4
rect 2730 -62 2784 0
rect 2914 -60 2968 2
rect 3110 -70 3164 -8
rect 3302 -66 3356 -4
rect 3494 -60 3548 2
rect 3686 -60 3740 2
rect 1862 -186 1914 -132
rect 2054 -182 2106 -128
rect 2244 -186 2296 -132
rect 2432 -190 2484 -136
rect 2628 -184 2680 -130
rect 2822 -188 2874 -134
rect 3014 -192 3066 -138
rect 3210 -188 3262 -134
rect 3402 -188 3454 -134
rect 3586 -188 3638 -134
rect 1496 -440 1568 -368
<< metal2 >>
rect 1500 1116 1572 1122
rect 1266 770 1346 776
rect 1266 350 1346 690
rect 1500 684 1572 1044
rect 1772 800 1828 810
rect 1964 804 2020 814
rect 1762 748 1772 800
rect 1828 748 1964 800
rect 1772 732 1828 742
rect 2150 806 2204 816
rect 2020 748 2150 800
rect 1964 736 2020 746
rect 2352 802 2406 812
rect 2204 748 2352 800
rect 2150 734 2204 744
rect 2540 802 2594 812
rect 2406 748 2540 800
rect 2352 730 2406 740
rect 2736 806 2790 816
rect 2594 748 2736 800
rect 2540 730 2594 740
rect 2920 808 2974 818
rect 2790 748 2920 800
rect 2736 734 2790 744
rect 3116 800 3170 808
rect 3308 802 3362 812
rect 2974 798 3308 800
rect 2974 748 3116 798
rect 2920 736 2974 746
rect 3170 748 3308 798
rect 3116 726 3170 736
rect 3500 808 3554 818
rect 3362 748 3500 800
rect 3308 730 3362 740
rect 3692 808 3746 818
rect 3554 748 3692 800
rect 3500 736 3554 746
rect 3746 748 4068 800
rect 3692 736 3746 746
rect 2060 684 2112 688
rect 2634 684 2686 686
rect 1500 678 3896 684
rect 1500 674 2060 678
rect 1500 620 1868 674
rect 1920 624 2060 674
rect 2112 676 3896 678
rect 2112 674 2634 676
rect 2112 624 2250 674
rect 1920 620 2250 624
rect 2302 670 2634 674
rect 2302 620 2438 670
rect 1500 616 2438 620
rect 2490 622 2634 670
rect 2686 672 3896 676
rect 2686 622 2828 672
rect 2490 618 2828 622
rect 2880 668 3216 672
rect 2880 618 3020 668
rect 2490 616 3020 618
rect 1500 614 3020 616
rect 3072 618 3216 668
rect 3268 618 3408 672
rect 3460 618 3592 672
rect 3644 618 3896 672
rect 3072 614 3896 618
rect 1500 612 3896 614
rect 1868 610 1920 612
rect 2250 610 2302 612
rect 2438 606 2490 612
rect 2828 608 2880 612
rect 3020 604 3072 612
rect 3216 608 3268 612
rect 3408 608 3460 612
rect 3592 608 3644 612
rect 4016 420 4068 748
rect 1266 270 1542 350
rect 1622 270 1628 350
rect 1266 -52 1346 270
rect 3994 227 4088 420
rect 3994 200 4119 227
rect 4016 110 4119 200
rect 1766 -6 1822 4
rect 1958 -2 2014 8
rect 1756 -58 1766 -6
rect 1822 -58 1958 -6
rect 1766 -74 1822 -64
rect 2144 0 2198 10
rect 2014 -58 2144 -6
rect 1958 -70 2014 -60
rect 2346 -4 2400 6
rect 2198 -58 2346 -6
rect 2144 -72 2198 -62
rect 2534 -4 2588 6
rect 2400 -58 2534 -6
rect 2346 -76 2400 -66
rect 2730 0 2784 10
rect 2588 -58 2730 -6
rect 2534 -76 2588 -66
rect 2914 2 2968 12
rect 2784 -58 2914 -6
rect 2730 -72 2784 -62
rect 3110 -6 3164 2
rect 3302 -4 3356 6
rect 2968 -8 3302 -6
rect 2968 -58 3110 -8
rect 2914 -70 2968 -60
rect 3164 -58 3302 -8
rect 3110 -80 3164 -70
rect 3494 2 3548 12
rect 3356 -58 3494 -6
rect 3302 -76 3356 -66
rect 3686 2 3740 12
rect 3548 -58 3686 -6
rect 3494 -70 3548 -60
rect 4006 -6 4119 110
rect 3740 -58 4119 -6
rect 3686 -70 3740 -60
rect 4006 -97 4119 -58
rect 4006 -102 4058 -97
rect 2054 -122 2106 -118
rect 2628 -122 2680 -120
rect 1266 -138 1346 -132
rect 1496 -128 3890 -122
rect 1496 -132 2054 -128
rect 1496 -186 1862 -132
rect 1914 -182 2054 -132
rect 2106 -130 3890 -128
rect 2106 -132 2628 -130
rect 2106 -182 2244 -132
rect 1914 -186 2244 -182
rect 2296 -136 2628 -132
rect 2296 -186 2432 -136
rect 1496 -190 2432 -186
rect 2484 -184 2628 -136
rect 2680 -134 3890 -130
rect 2680 -184 2822 -134
rect 2484 -188 2822 -184
rect 2874 -138 3210 -134
rect 2874 -188 3014 -138
rect 2484 -190 3014 -188
rect 1496 -192 3014 -190
rect 3066 -188 3210 -138
rect 3262 -188 3402 -134
rect 3454 -188 3586 -134
rect 3638 -188 3890 -134
rect 3066 -192 3890 -188
rect 1496 -194 3890 -192
rect 1496 -368 1568 -194
rect 1862 -196 1914 -194
rect 2244 -196 2296 -194
rect 2432 -200 2484 -194
rect 2822 -198 2874 -194
rect 3014 -202 3066 -194
rect 3210 -198 3262 -194
rect 3402 -198 3454 -194
rect 3586 -198 3638 -194
rect 1496 -446 1568 -440
use sky130_fd_pr__pfet_01v8_8DVCWJ  sky130_fd_pr__pfet_01v8_8DVCWJ_0
timestamp 1711967491
transform 1 0 2757 0 1 707
box -1127 -319 1127 319
use sky130_fd_pr__nfet_01v8_YTLFGX  XM2
timestamp 1711967491
transform 1 0 2751 0 1 -100
box -1127 -310 1127 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM3
timestamp 1711967491
transform 1 0 987 0 1 717
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM4
timestamp 1711967491
transform 1 0 983 0 1 -92
box -211 -310 211 310
<< labels >>
flabel metal1 -138 -768 62 -568 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 76 192 276 392 0 FreeSans 256 0 0 0 IN
port 3 nsew
flabel metal1 4142 240 4342 440 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 -134 1208 66 1408 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal2 1266 -52 1346 690 0 FreeSans 320 0 0 0 not_in
<< end >>
