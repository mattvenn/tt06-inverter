magic
tech sky130A
magscale 1 2
timestamp 1712075644
<< metal1 >>
rect 18568 6436 18868 6442
rect 18868 6432 19868 6436
rect 18868 6140 19870 6432
rect 18868 6136 19868 6140
rect 18568 6130 18868 6136
rect 19710 5186 20008 5406
rect 23862 5302 24240 5422
rect 19710 5138 19778 5186
rect 19772 5066 19778 5138
rect 19898 5138 20008 5186
rect 24120 5254 24240 5302
rect 26896 5254 27016 5260
rect 19898 5066 19904 5138
rect 24120 5134 26896 5254
rect 26896 5128 27016 5134
rect 19220 4236 19872 4458
rect 18936 4230 19872 4236
rect 19236 4158 19872 4230
rect 19236 3930 19520 4158
rect 18936 3924 19236 3930
<< via1 >>
rect 18568 6136 18868 6436
rect 19778 5066 19898 5186
rect 26896 5134 27016 5254
rect 18936 3930 19236 4230
<< metal2 >>
rect 17919 6436 18209 6440
rect 17914 6431 18568 6436
rect 17914 6141 17919 6431
rect 18209 6141 18568 6431
rect 17914 6136 18568 6141
rect 18868 6136 18874 6436
rect 17919 6132 18209 6136
rect 19778 5186 19898 5192
rect 26890 5134 26896 5254
rect 27016 5134 27022 5254
rect 19778 5035 19898 5066
rect 19774 4925 19783 5035
rect 19893 4925 19902 5035
rect 19778 4920 19898 4925
rect 26896 4249 27016 5134
rect 18675 4230 18965 4234
rect 18670 4225 18936 4230
rect 18670 3935 18675 4225
rect 18670 3930 18936 3935
rect 19236 3930 19242 4230
rect 26892 4139 26901 4249
rect 27011 4139 27020 4249
rect 26896 4134 27016 4139
rect 18675 3926 18965 3930
<< via2 >>
rect 17919 6141 18209 6431
rect 19783 4925 19893 5035
rect 18675 3935 18936 4225
rect 18936 3935 18965 4225
rect 26901 4139 27011 4249
<< metal3 >>
rect 6563 6436 6861 6441
rect 6562 6435 18214 6436
rect 6562 6137 6563 6435
rect 6861 6431 18214 6435
rect 6861 6141 17919 6431
rect 18209 6141 18214 6431
rect 6861 6137 18214 6141
rect 6562 6136 18214 6137
rect 6563 6131 6861 6136
rect 19778 5035 19898 5040
rect 19778 4925 19783 5035
rect 19893 4925 19898 5035
rect 19778 4793 19898 4925
rect 19773 4675 19779 4793
rect 19897 4675 19903 4793
rect 19778 4674 19898 4675
rect 26896 4249 27016 4254
rect 18393 4230 18691 4235
rect 18392 4229 18970 4230
rect 18392 3931 18393 4229
rect 18691 4225 18970 4229
rect 18965 3935 18970 4225
rect 18691 3931 18970 3935
rect 18392 3930 18970 3931
rect 26896 4139 26901 4249
rect 27011 4139 27016 4249
rect 18393 3925 18691 3930
rect 26896 1705 27016 4139
rect 26891 1587 26897 1705
rect 27015 1587 27021 1705
rect 26896 1586 27016 1587
<< via3 >>
rect 6563 6137 6861 6435
rect 19779 4675 19897 4793
rect 18393 4225 18691 4229
rect 18393 3935 18675 4225
rect 18675 3935 18691 4225
rect 18393 3931 18691 3935
rect 26897 1587 27015 1705
<< metal4 >>
rect 798 44660 858 45152
rect 1534 44660 1594 45152
rect 2270 44660 2330 45152
rect 3006 44660 3066 45152
rect 3742 44660 3802 45152
rect 4478 44660 4538 45152
rect 5214 44660 5274 45152
rect 5950 44660 6010 45152
rect 6686 44660 6746 45152
rect 7422 44660 7482 45152
rect 8158 44660 8218 45152
rect 8894 44660 8954 45152
rect 9630 44660 9690 45152
rect 10366 44660 10426 45152
rect 11102 44660 11162 45152
rect 11838 44660 11898 45152
rect 12574 44660 12634 45152
rect 13310 44660 13370 45152
rect 14046 44660 14106 45152
rect 14782 44660 14842 45152
rect 15518 44660 15578 45152
rect 16254 44660 16314 45152
rect 16990 44660 17050 45152
rect 17726 44660 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 742 44284 17786 44660
rect 200 6436 500 44152
rect 200 6435 6862 6436
rect 200 6137 6563 6435
rect 6861 6137 6862 6435
rect 200 6136 6862 6137
rect 200 1000 500 6136
rect 9800 4230 10100 44284
rect 17726 44270 17786 44284
rect 19778 4793 19898 4794
rect 19778 4675 19779 4793
rect 19897 4675 19898 4793
rect 9800 4229 18692 4230
rect 9800 3931 18393 4229
rect 18691 3931 18692 4229
rect 9800 3930 18692 3931
rect 9800 1000 10100 3930
rect 19778 3206 19898 4675
rect 19778 3086 31432 3206
rect 26896 1705 27016 1706
rect 26896 1587 26897 1705
rect 27015 1587 27016 1705
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 1587
rect 31312 0 31432 3086
use inverter  inverter_0
timestamp 1712074259
transform 1 0 19706 0 1 4996
box -236 -828 4448 1468
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
