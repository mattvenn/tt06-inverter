magic
tech sky130A
magscale 1 2
timestamp 1712322988
<< error_p >>
rect -29 181 29 187
rect -29 147 -17 181
rect -29 141 29 147
rect -29 -147 29 -141
rect -29 -181 -17 -147
rect -29 -187 29 -181
<< nwell >>
rect -213 -319 213 319
<< pmos >>
rect -17 -100 17 100
<< pdiff >>
rect -75 88 -17 100
rect -75 -88 -63 88
rect -29 -88 -17 88
rect -75 -100 -17 -88
rect 17 88 75 100
rect 17 -88 29 88
rect 63 -88 75 88
rect 17 -100 75 -88
<< pdiffc >>
rect -63 -88 -29 88
rect 29 -88 63 88
<< nsubdiff >>
rect -177 249 -81 283
rect 81 249 177 283
rect -177 187 -143 249
rect 143 187 177 249
rect -177 -249 -143 -187
rect 143 -249 177 -187
rect -177 -283 -81 -249
rect 81 -283 177 -249
<< nsubdiffcont >>
rect -81 249 81 283
rect -177 -187 -143 187
rect 143 -187 177 187
rect -81 -283 81 -249
<< poly >>
rect -33 181 33 197
rect -33 147 -17 181
rect 17 147 33 181
rect -33 131 33 147
rect -17 100 17 131
rect -17 -131 17 -100
rect -33 -147 33 -131
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect -33 -197 33 -181
<< polycont >>
rect -17 147 17 181
rect -17 -181 17 -147
<< locali >>
rect -177 249 -81 283
rect 81 249 177 283
rect -177 187 -143 249
rect 143 187 177 249
rect -33 147 -17 181
rect 17 147 33 181
rect -63 88 -29 104
rect -63 -104 -29 -88
rect 29 88 63 104
rect 29 -104 63 -88
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect -177 -249 -143 -187
rect 143 -249 177 -187
rect -177 -283 -81 -249
rect 81 -283 177 -249
<< viali >>
rect -17 147 17 181
rect -63 -88 -29 88
rect 29 -88 63 88
rect -17 -181 17 -147
<< metal1 >>
rect -29 181 29 187
rect -29 147 -17 181
rect 17 147 29 181
rect -29 141 29 147
rect -69 88 -23 100
rect -69 -88 -63 88
rect -29 -88 -23 88
rect -69 -100 -23 -88
rect 23 88 69 100
rect 23 -88 29 88
rect 63 -88 69 88
rect 23 -100 69 -88
rect -29 -147 29 -141
rect -29 -181 -17 -147
rect 17 -181 29 -147
rect -29 -187 29 -181
<< properties >>
string FIXED_BBOX -160 -266 160 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.17 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
